    function new(string name, uvm_component parent);
      super.new(name, parent);
    endfunction : new
