class component extends uvm_component;
    `uvm_component_utils(component)

    function new(string name, uvm_component parent);
      super.new(name, parent);
    endfunction : new


endclass : component
